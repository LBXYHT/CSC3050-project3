`timescale 1ns/1ps

module alu_test;

reg [31:0] instruction, reg1, reg2;

wire [31:0] final_result;
wire [2:0] flag; 
//wire zero;
//wire overflow;
//wire neg;

ALU testalu(instruction, reg1, reg2, final_result, flag);

initial
begin

$display("instruction: reg1: reg2: final_result: flag");
$monitor("%h:%h:%h:%b:%b",instruction, reg1, reg2, final_result, flag);

//add1
#10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0000;
reg1<=32'b1000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b1011_1111_1111_1111_1111_1111_1111_1110;

//add2
#10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0000;
reg1<=32'b0100_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b0111_1111_1111_1111_1111_1111_1111_1110;

//add3
#10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0000;
reg1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b1000_1111_1111_1111_1111_1111_1111_1110;

//addu
#10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0001;
reg1<=32'b1000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b1011_1111_1111_1111_1111_1111_1111_1110;

//and
#10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0100;
reg1<=32'b0000_0000_1111_0000_0000_1111_0000_1010;
reg2<=32'b1011_1111_1111_1111_1111_1111_1111_1110;

//nor
#10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0111;
reg1<=32'b1000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b1011_1111_1111_1111_1111_1111_1111_1110;

//or
#10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0101;
reg1<=32'b1000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b1011_0000_1111_1111_1111_0000_1111_1110;

//sll1
#10 instruction<=32'b0000_0000_0010_0001_0000_0000_1100_0000;
reg1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b1011_0000_0000_1111_0000_0000_0001_1000;

//sll2
#10 instruction<=32'b0000_0000_0000_0000_0000_0000_1100_0000;
reg1<=32'b0110_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b0000_0000_0000_0000_0000_0000_0001_1000;

//sllv
#10 instruction<=32'b0000_0000_0010_0001_0000_0000_0000_0100;
reg1<=32'b0000_0000_0000_0000_0000_0000_0000_1110;
reg2<=32'b1011_0111_1001_0000_1111_1111_1000_0000;

//slt1
#10 instruction<=32'b0000_0000_0000_0000_0000_0000_0010_1010;
reg1<=32'b1100_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b1011_1111_1111_1111_1111_1111_1111_1110;

//slt2
#10 instruction<=32'b0000_0000_0010_0000_0000_0000_0010_1010;
reg1<=32'b1000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b0011_1111_1111_1111_1111_1111_1111_1110;

//sltu1
#10 instruction<=32'b0000_0000_0000_0000_0000_0000_0010_1011;
reg1<=32'b1000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b0000_0000_0000_0000_0000_0000_0000_0010;

//sltu2
#10 instruction<=32'b0000_0000_0010_0000_0000_0000_0010_1011;
reg1<=32'b0000_0000_0000_0000_0000_0000_0000_0110;
reg2<=32'b0000_0000_0000_0000_0000_0000_0000_0010;

//sra
#10 instruction<=32'b0000_0000_0000_0001_0000_0000_1000_0011;
reg1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b0011_1111_1111_1111_1111_1111_1111_1110;

//srav
#10 instruction<=32'b0000_0000_0000_0001_0000_0010_0000_0111;
reg1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b0011_1111_1111_1111_1111_1111_1111_1110;

//srl1
#10 instruction<=32'b0000_0000_0000_0001_0000_0000_0000_0010;
reg1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b0011_1111_1111_1111_1111_1111_1111_1110;

//srl2
#10 instruction<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
reg1<=32'b1111_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b0000_0000_0000_0000_0000_0000_0011_0011;

//srlv
#10 instruction<=32'b0000_0000_0000_0001_0000_0000_0000_0110;
reg1<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
reg2<=32'b0011_1111_1111_1111_1111_1111_1111_1110;

//sub1
#10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0010;
reg1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//sub2
#10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0010;
reg1<=32'b1000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b0000_0000_0000_0011_1100_1100_0000_1110;

//sub3
#10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0010;
reg1<=32'b0111_1111_1111_1110_0000_0000_0000_0010;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//subu
#10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0011;
reg1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//xor
#10 instruction<=32'b0000_0000_0000_0000_0000_0000_0010_0110;
reg1<=32'b0000_0000_0000_0000_0011_0000_0000_0010;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//addi1
#10 instruction<=32'b0010_0000_0000_0000_0000_0000_0010_0010;
reg1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//addi2
#10 instruction<=32'b0010_0000_0000_0000_1111_1111_0010_0010;
reg1<=32'b1000_0000_0000_0000_0000_0000_0100_0010;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//addi3
#10 instruction<=32'b0010_0000_0010_0000_0111_0000_0010_0010;
reg1<=32'b1000_0000_0000_0011_1100_1100_0000_1110;
reg2<=32'b0111_1111_1111_1111_1111_1111_0000_0010;

//addiu
#10 instruction<=32'b0010_0100_0000_0001_1000_0000_0010_0010;
reg1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//andi
#10 instruction<=32'b0011_0000_0000_0000_1111_0010_0010_0110;
reg1<=32'b0000_0000_0000_0000_1110_1100_0110_0110;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//beq1
#10 instruction<=32'b0001_0000_0000_0000_0000_0000_0010_0010;
reg1<=32'b1000_0000_0011_0111_0110_0000_0000_0010;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//beq2
#10 instruction<=32'b0001_0000_0000_0000_0000_0000_0010_0010;
reg1<=32'b1000_0000_0011_0111_0110_0000_0000_0010;
reg2<=32'b1000_0000_0011_0111_0110_0000_0000_0010;

//bne1
#10 instruction<=32'b0001_0100_0000_0000_0000_0000_0010_0010;
reg1<=32'b1000_0000_0011_0111_0110_0000_0000_0010;
reg2<=32'b1000_0000_0011_0111_0110_0000_0000_0010;

//bne2
#10 instruction<=32'b0001_0100_0000_0000_0000_0000_0010_0010;
reg1<=32'b0000_1000_0011_0111_0110_0000_0000_0010;
reg2<=32'b1000_0010_0011_0101_1100_1100_0000_1111;

//lw
#10 instruction<=32'b1000_1100_0000_0000_0000_0000_0010_0010;
reg1<=32'b1000_0000_0011_0111_0110_0000_0000_0010;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//ori
#10 instruction<=32'b0011_0100_0000_0000_0000_0000_0010_0010;
reg1<=32'b1000_0000_0011_0111_0110_0000_0000_0010;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//slti1
#10 instruction<=32'b0010_1000_0000_0000_0000_0000_0010_0010;
reg1<=32'b0000_0000_0011_0111_0110_0000_0010_0010;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//slti2
#10 instruction<=32'b0010_1000_0010_0000_0000_0000_0010_0010;
reg1<=32'b0000_0000_0011_0111_0110_0000_0010_0010;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//sltiu1
#10 instruction<=32'b0010_1100_0000_0000_1000_0000_0010_0010;
reg1<=32'b0000_0000_0011_0111_0110_0000_0010_0010;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//sltiu2
#10 instruction<=32'b0010_1100_0010_0000_0000_0000_0010_0010;
reg1<=32'b0000_0000_0011_0111_0110_0000_0010_0010;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//sw
#10 instruction<=32'b1010_1100_0000_0000_0000_0000_0010_0010;
reg1<=32'b0000_0000_0011_0111_0110_0000_0010_0010;
reg2<=32'b1000_0000_0000_0011_1100_1100_0000_1110;

//xori
#10 instruction<=32'b0011_1000_0000_0000_0000_0000_0010_0010;
reg1<=32'b0000_0000_0011_0111_0110_0000_0010_0010;
reg2<=32'b1000_0000_0110_0000_0001_1100_0000_0110;



/*
#10 instruction<=32'b0000_0000_0000_0001_0001_0000_0100_0000;
gr1<=32'b0100_0000_0100_0000_0100_0000_0100_0000;

#10 instruction<=32'b0000_0000_0000_0001_0001_0001_0000_0000;
gr1<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
*/

#10 $finish;
end
endmodule